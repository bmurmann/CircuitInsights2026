.param id = 3.76e-04
.param w = 6.23e-05
.param l = 1.30e-07
.param nf = 13.0
.param rd = 1.00e+03
.param rs = 1.00e+04
.param cl = 2.00e-13
